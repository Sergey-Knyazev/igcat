REGIONS:	errors	(signed	/ unsigned)	(signed	/ unsigned)
FR1 start:	2	(-0.009	/ 0.009)	(-1.500	/ 1.500)
FR1 end:	1	(0.003	/ 0.003)	(1.000	/ 1.000)
CDR1 start:	1	(0.003	/ 0.003)	(1.000	/ 1.000)
CDR1 end:	0	(0.000	/ 0.000)	(0.000	/ 0.000)
FR2 start:	0	(0.000	/ 0.000)	(0.000	/ 0.000)
FR2 end:	0	(0.000	/ 0.000)	(0.000	/ 0.000)
CDR2 start:	0	(0.000	/ 0.000)	(0.000	/ 0.000)
CDR2 end:	2	(0.006	/ 0.006)	(1.000	/ 1.000)
FR3 start:	0	(0.000	/ 0.000)	(0.000	/ 0.000)
FR3 end:	24	(-0.003	/ 0.098)	(-0.042	/ 1.375)
CDR3 start:	29	(-0.006	/ 0.107)	(-0.069	/ 1.241)
CDR3 end:	0	(0.000	/ 0.000)	(0.000	/ 0.000)
FR4 start:	0	(0.000	/ 0.000)	(0.000	/ 0.000)
FR4 end:	39	(0.116	/ 0.116)	(1.000	/ 1.000)
